LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Processador IS
    PORT ( 
	        CLK : IN STD_LOGIC;
           RESET : IN STD_LOGIC;
           FUNCTION_CODE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
           DATA_IN : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
           DATA_OUT : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
			  
			 );
			 
END Processador;

ARCHITECTURE BEHAVIORAL OF Processador IS

    SIGNAL R1, R2, R3, A, G: STD_LOGIC_VECTOR (3 DOWNTO 0);
    SIGNAL LOAD_R1, LOAD_R2, LOAD_R3, LOAD_A, LOAD_G, ADD_SUB, SWAP_START : STD_LOGIC;
    SIGNAL ULA_OUT : STD_LOGIC_VECTOR (3 DOWNTO 0);
    SIGNAL ULA_CARRY : STD_LOGIC;

    COMPONENT REGISTRADOR
	 
        PORT ( 
		         CLK, LOAD : IN STD_LOGIC;
					RESET : in STD_LOGIC;
					D : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
					Q : OUT STD_LOGIC_VECTOR (3 DOWNTO 0) 
				  );
				  
    END COMPONENT;

    COMPONENT ULA
	 
        PORT ( 
					A: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
               B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
               ADD_SUB : IN STD_LOGIC;
               F: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
					CARRY_OUT: OUT STD_LOGIC
				  );
				  
    END COMPONENT;

    COMPONENT UnidadeDeControle IS

    PORT ( 
           CLK : IN STD_LOGIC;
			  RESET : IN STD_LOGIC;
           FUNCTION_CODE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
           LOAD_R1 : OUT STD_LOGIC;
           LOAD_R2 : OUT STD_LOGIC;
           LOAD_R3 : OUT STD_LOGIC;
			  LOAD_A  : OUT STD_LOGIC;
			  LOAD_G  : OUT STD_LOGIC;
           ADD_SUB : OUT STD_LOGIC;
			  SWAP_START : OUT STD_LOGIC
         );
			
	 END COMPONENT UnidadeDeControle;
	 
	 COMPONENT SWAP IS
    PORT (
        CLOCK : IN STD_LOGIC;
        RESET : IN STD_LOGIC;
        START : IN STD_LOGIC;
        R1_IN : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
        R2_IN : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
        R1_OUT : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
        R2_OUT : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
        
       );
	 END COMPONENT SWAP;


BEGIN

    -- INSTANCIAÇÃO DOS REGISTRADORES
	 
    REG1 : REGISTRADOR PORT MAP(CLK, LOAD_R1, RESET, DATA_IN, R1);
    REG2 : REGISTRADOR PORT MAP(CLK, LOAD_R2, RESET, DATA_IN, R2);
    REG3 : REGISTRADOR PORT MAP(CLK, LOAD_R3, RESET, DATA_IN, R3);
	 RegA : REGISTRADOR port map(CLK, LOAD_A , RESET, R2     ,  A); 
    RegG : REGISTRADOR port map(CLK, LOAD_G , RESET, ULA_OUT,  G); 

    -- INSTANCIAÇÃO DA ULA
	 
    ULA0 : ULA PORT MAP(A, R1, ADD_SUB, ULA_OUT, ULA_CARRY);

    -- SWAP
	 
	 -- Instanciação do SWAP
    SWAP0 : SWAP PORT MAP(CLK, RESET, SWAP_START, R1, R2);  -- FALTA DEFINIR AS SAÍDAS DO SWAP E ATUALIZAR O VALOR DE R1 E R2
	 
    
    -- INSTANCIAÇÃO DA UNIDADE DE CONTROLE
    CONTROL_UNIT : UnidadeDeControle PORT MAP(CLK, RESET, FUNCTION_CODE, LOAD_R1, LOAD_R2, LOAD_R3, LOAD_A, LOAD_G, ADD_SUB, SWAP_START);

    -- SAÍDA DE DADOS
	 
    DATA_OUT <= G;
	 
END BEHAVIORAL;
